`ifndef BRCTYPE
    localparam BEQ  = 3'b000;
    localparam BNE  = 3'b001;
    localparam BLT  = 3'b100;
    localparam BGE  = 3'b101;
    localparam BLTU = 3'b110;
    localparam BGEU = 3'b111;
    localparam BNONE = 3'b010;
`define BRCTYPE
`endif
