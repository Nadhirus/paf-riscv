`ifndef ALUTYPE
localparam ADD = 4'b0000;
localparam SUB = 4'b1000;
localparam SLL = 4'b0001;
localparam SLT = 4'b0010;
localparam SLTU= 4'b0011;
localparam XOR = 4'b0100;
localparam SRL = 4'b0101;
localparam SRA = 4'b1101;
localparam  OR = 4'b0110;
localparam AND = 4'b0111;
`define ALUTYPE
`endif
